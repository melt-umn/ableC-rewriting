grammar edu:umn:cs:melt:exts:ableC:rewriting;

exports edu:umn:cs:melt:exts:ableC:rewriting:concretesyntax;
exports edu:umn:cs:melt:exts:ableC:rewriting:abstractsyntax;

exports edu:umn:cs:melt:exts:ableC:templating;
exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes;
exports edu:umn:cs:melt:exts:ableC:closure;
